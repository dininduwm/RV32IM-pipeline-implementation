`timescale 1ns/100ps

module branch_select(DATA1, DATA2, SELECT, MUX_OUT);

    input [31:0] DATA1, DATA2;
    input [3:0] SELECT;
    output reg MUX_OUT;

    // TODO: implement the function



endmodule