`timescale 1ns/100ps

module adder(INPUT1, INPUT2, RESULT); // adder module

    input [31:0] INPUT1, INPUT2; // declare inputs
    output reg [31:0] RESULT;    // declare outputs

    always @(*) 
    begin
      // TODO : set the time delay
      #2 RESULT = INPUT1 + INPUT2; // add two numbers 
    end

endmodule