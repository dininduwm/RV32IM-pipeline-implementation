`timescale 1ns/100ps

module twosComp(INPUT, RESULT); //change this
    input [31:0] INPUT;       //declare inputs
    output reg [31:0] RESULT; //declare outputs

    always @ (INPUT)
    begin
      // TODO : set the time delay
      #1 RESULT = ~INPUT + 1; // 2s comp negative
    end

endmodule